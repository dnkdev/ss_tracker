module main

// import web
// import database
// import parser
import bot

fn main() {
	bot.start_bot()!
	// user := User{telegram_id: 100, lang: .en}
	// users := get_users(db)!
	// println(user_exist(db,user))
	// add_user(db,user)
	// println(users)

	// web.start_server(web.new_app())

	// mut result := get_category()
	// url := 'https://ss.com${result}'
	// println(url)
	// mut response := http.get(url) !
	// //result := http.get('https://ss.com') or{panic(err)}
	// mut file := os.open_file('result.html','w') !
	// defer{
	// 	file.close()
	// }
	// file.write_string(response.body) !
	// //tbot.main()
}
