module main

fn main() {
	start_bot() or {
		panic(err)
	}
}
