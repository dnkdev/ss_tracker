module main

import bot

fn main() {
	bot.start_bot()!
}
